`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/07/2024 12:00:57 PM
// Design Name: 
// Module Name: object
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module object #( 

// Image resolution
parameter HRES = 1280,
parameter VRES = 720,

// Object Color
parameter COLOR = 24'h 00FF90,

// Paddle Height
parameter PADDLE_H = 20
)
(
    input pixel_clk,
    input rst,
    input fsync, 
    
    // Paddle location
    input signed [11:0] hpos, 
    input signed [11:0] vpos, 
    input [1:0] random_number, // Input port for the random number generated by LFSR

    output [7:0] pixel [0:2], 
    
    output [11:0] left_edge,

    
    output active, 
    
    input player_1_score
    
);
    localparam OBJ_SIZE = 50; 
    localparam [1:0] DOWN_RIGHT = 2'b00; 
    localparam [1:0] DOWN_LEFT  = 2'b01; 
    localparam [1:0] UP_RIGHT   = 2'b10; 
    localparam [1:0] UP_LEFT    = 2'b11;
    
    // Velocity of ball, 12 pixels per clock cycle
    localparam VEL = 8; 
    
    // Paddle location in horizontal/vertical format
    reg signed [11 : 0  ] lhpos; // left horizontal position 
    reg signed [11 : 0  ] rhpos; // right horizonat position 
    reg signed [11 : 0  ] tvpos; // top vertical position 
    reg signed [11 : 0  ] bvpos; // bottom vertical position
    
    
    reg [1 : 0 ] dir ; // direction of object 

    
   
    always @(posedge pixel_clk)     
//begin if(vpos <= PADDLE_H -40 && active)
//    begin
//case (random_number)
//        // Case 1: Active and random_number = 2'b01
//        2'b00: begin
//            lhpos = 100;
//            rhpos = 100 + OBJ_SIZE - 1;
//            tvpos = 100;
//            bvpos = 100 + OBJ_SIZE - 1;
//            dir = DOWN_RIGHT;
//        end
//        // Case 2: Active and random_number = 2'b00
//        2'b01: begin
//            lhpos = 1000;
//            rhpos = 1000 + OBJ_SIZE - 1;
//            tvpos = 220;
//            bvpos = 220 + OBJ_SIZE - 1;
//            dir = DOWN_LEFT;
//        end
//        // Case 3: Active and random_number = 2'b10
//        2'b10: begin
//            lhpos = 500;
//            rhpos = 500 + OBJ_SIZE - 1;
//            tvpos = 580;
//            bvpos = 580 + OBJ_SIZE - 1;
//            dir = UP_RIGHT;
//        end
//        // Case 4: Active and random_number = 2'b11
//        2'b11: begin
//            lhpos = 600;
//            rhpos = 600 + OBJ_SIZE - 1;
//            tvpos = 580;
//            bvpos = 580 + OBJ_SIZE - 1;
//            dir = UP_RIGHT;
//        end
//        // Default case: Inactive
//        default: begin
//            // Do nothing when not active
//        end
//    endcase
//    end
begin
    if(player_1_score) begin 
        // Generate a random number between 1 and 3 inclusive
        // Set values based on the random number
        case(random_number)
            2'b01: begin
                lhpos <= 100;
                rhpos <= 100 + OBJ_SIZE - 1;
                tvpos <= 100;
                bvpos <= 100 + OBJ_SIZE - 1;
                dir   <= DOWN_RIGHT;       // Reset direction to DOWN_RIGHT
            end
            2'b00: begin
                lhpos <= 1000;
                rhpos <= 1000 + OBJ_SIZE - 1;
                tvpos <= 220;
                bvpos <= 220 + OBJ_SIZE - 1;
                dir   <= DOWN_LEFT;       // Reset direction to DOWN_LEFT
            end
            2'b10: begin
                lhpos <= 500;
                rhpos <= 500 + OBJ_SIZE - 1;
                tvpos <= 580;
                bvpos <= 580 + OBJ_SIZE - 1;
                dir   <= UP_RIGHT;       // Reset direction to UP_RIGHT
            end
            2'b11: begin
                lhpos <= 600;
                rhpos <= 600 + OBJ_SIZE - 1;
                tvpos <= 580;
                bvpos <= 580 + OBJ_SIZE - 1;
                dir   <= UP_RIGHT;       // Reset direction to UP_RIGHT
            end
            default: begin
                // Default case (should not happen)
                lhpos <= 1000;
                rhpos <= 1000 + OBJ_SIZE - 1;
                tvpos <= 1000;
                bvpos <= 1000 + OBJ_SIZE - 1;
                dir   <= DOWN_RIGHT;       // Reset direction to DOWN_RIGHT
            end
        endcase
    end else if (fsync) begin 
             if(dir == DOWN_RIGHT) begin 
                if (bvpos == VRES - PADDLE_H) begin 
                    dir <= UP_RIGHT; 
                end else if (rhpos == HRES - 1) begin 
                    dir <= DOWN_LEFT;
                end 
            end 

            // Down Left
            else if(dir == DOWN_LEFT) begin 
                if (bvpos == VRES - PADDLE_H) begin 
                    dir <= UP_LEFT; 
                end else if (lhpos == 0) begin 
                    dir <= DOWN_RIGHT;
                end 
            end 

            // Top Right FOR BOTH TOP POSITIONS NEED TO MAKE SURE IT DOESN"T BOUNCE OFF THE TOP
            else if(dir == UP_RIGHT) begin 
                if (tvpos == 0) begin 
                    dir <= DOWN_RIGHT; 
                end else if (rhpos == HRES - 1) begin 
                    dir <= UP_LEFT;
                end 
            end 

            // Top left
            else if(dir == UP_LEFT) begin 
                if (tvpos == 0) begin 
                    dir <= DOWN_LEFT; 
                end else if (lhpos == 0) begin 
                    dir <= UP_RIGHT;
                end 
            end

 
            // Example Code
            if  (dir == DOWN_RIGHT) begin // Check if new ball location is still within bounds 
                if ( ( rhpos + VEL) <= HRES  - 1 && (bvpos + VEL) <= VRES - PADDLE_H) begin 
                    lhpos <= lhpos + VEL ; 
                    rhpos <= rhpos + VEL ; 
                    tvpos <= tvpos + VEL ; 
                    bvpos <= bvpos + VEL ; 
                
                //end else if (...) begin 
                //end else if
               end  else if ( ( rhpos + VEL) > HRES  - 1) begin
                    lhpos <= HRES -OBJ_SIZE ; 
                    rhpos <= HRES - 1 ; 
                    tvpos <= tvpos + VEL ; 
                    bvpos <= bvpos + VEL ;
               // ....
            end else if ((bvpos + VEL) > VRES - PADDLE_H) begin
                    lhpos <= lhpos + VEL; 
                    rhpos <= rhpos + VEL; 
                    tvpos <= VRES - PADDLE_H - OBJ_SIZE + 1; 
                    bvpos <= VRES - PADDLE_H; 
            end 
            end

            else if (dir == UP_RIGHT) begin
                if ((rhpos + VEL) <= HRES - 1 && (tvpos - VEL) >= 0) begin
                    lhpos <= lhpos + VEL ; 
                    rhpos <= rhpos + VEL ; 
                    tvpos <= tvpos - VEL ; 
                    bvpos <= bvpos - VEL ; 
                end else if ((rhpos + VEL) > HRES-1 ) begin
                    lhpos <= HRES -OBJ_SIZE ; 
                    rhpos <= HRES - 1 ; 
                    tvpos <= tvpos - VEL ; 
                    bvpos <= bvpos - VEL ;
                end else if ((tvpos - VEL) <0 ) begin  
                    tvpos <= 0;
                    bvpos <= OBJ_SIZE -1 ;
                    lhpos <= lhpos + VEL; 
                    rhpos <= rhpos + VEL; 
               end
               end
            
            else if (dir == UP_LEFT) begin
                if ((lhpos - VEL) >= 0 && (tvpos - VEL) >= 0) begin
                    lhpos <= lhpos - VEL ; 
                    rhpos <= rhpos - VEL ; 
                    tvpos <= tvpos - VEL ; 
                    bvpos <= bvpos - VEL ; 
                end  else if ((lhpos - VEL) <0 ) begin  
                    lhpos <= 0;
                    rhpos <= OBJ_SIZE -1 ;
                    tvpos <= tvpos - VEL; 
                    bvpos <= bvpos - VEL; 
                end  else if ((tvpos - VEL) <0 ) begin  
                    tvpos <= 0;
                    bvpos <= OBJ_SIZE -1 ;
                    lhpos <= lhpos - VEL; 
                    rhpos <= rhpos - VEL; 
            end 
            

            end else if (dir == DOWN_LEFT) begin
                if ((lhpos - VEL) >= 0 && (bvpos + VEL) <= VRES - PADDLE_H) begin
                    lhpos <= lhpos - VEL ; 
                    rhpos <= rhpos - VEL ; 
                    tvpos <= tvpos + VEL ; 
                    bvpos <= bvpos + VEL ; 
                end else if ((lhpos - VEL) <0 ) begin  
                    lhpos <= 0;
                    rhpos <= OBJ_SIZE -1 ;
                    tvpos <= tvpos + VEL; 
                    bvpos <= bvpos + VEL; 
                end else if ((bvpos + VEL) > VRES - PADDLE_H) begin
                    lhpos <= lhpos - VEL; 
                    rhpos <= rhpos - VEL; 
                    tvpos <= VRES - PADDLE_H - OBJ_SIZE + 1; 
                    bvpos <= VRES - PADDLE_H; 

            end

          end 
        end 
    end 
    
                                 
    /* Active calculates whether the current pixel being updated by the HDMI controller is within the bounds of the ball's */
    /* Simple Example: If the ball is located at position 0,0 and vpos and rpos = 0, active will be high, placing a green pixel */
    assign active = (hpos >= lhpos && hpos <= rhpos && vpos >= tvpos && vpos <= bvpos ) ? 1'b1 : 1'b0 ; 
    assign left_edge = lhpos;

    /* If active is high, set the RGB values for neon green */
    assign pixel [ 2 ] = (active) ? COLOR [ 23 : 16 ] : 8 'h00; //red 
    assign pixel [ 1 ] = (active) ? COLOR [ 15 : 8 ] : 8 'h00; //green 
    assign pixel [ 0 ] = (active) ? COLOR [ 7 : 0 ] : 8 'h00; //blue 
    
     
    
endmodule
